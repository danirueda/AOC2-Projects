----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:38:18 05/15/2014 
-- Design Name: 
-- Module Name:    UC_DMA - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity UC_DMA is
     Port ( clk : in  STD_LOGIC;
          reset : in  STD_LOGIC;
          empezar: in  STD_LOGIC;
          fin: in  STD_LOGIC; --
          L_E: in  STD_LOGIC;  -- 0 lectura de memoria, 1 escritura en memoria
          Bus_Req: in std_logic;        -- solicitud del mips
		  IO_sync: in std_logic; -- se�al de sincro con el perif�rico
		  update_done :out std_logic; --para actualizar el bit done al terminar una transferencia
		  DMA_send_data: out std_logic; -- env�o de los datos al bus
		  DMA_send_addr: out std_logic; -- env�o de la direcci�n al bus
		  DMA_Burst: out std_logic; -- se�al de modo r�faga la activa si le piden que transfiera m�s de 1 palabra
		  DMA_wait: out std_logic; -- se�al de espera para la MD
		  reset_count: out std_logic; -- pone el contador a 0
		  count_enable: out std_logic; -- incrementa el contador 
		  load_data: out std_logic; -- carga una plabara de memoria o de IO
		  DMA_MD_RE: out std_logic; -- enable lectura mem
		  DMA_MD_WE: out std_logic; -- enable escritura mem
		  DMA_IO_RE: out std_logic; -- enable lectura IO
		  DMA_IO_WE: out std_logic; -- enable escritura IO
		  DMA_sync: out std_logic -- se�al de sincro con el perif�rico
		  );
end UC_DMA;

architecture Behavioral of UC_DMA is
   --Si pon�is en el siguiente tipo el nombre de vuestros estados, los pod�is usar despu�s. Os pongo un ejemplo con algunos nombres. Cambiadlos, y a�adid los que necesit�is.
   type state_type is (INI, Escribir_IO, Leer_IO) ; 
   signal state, next_state : state_type; 
   
begin
 
 
-- registro de estado (en cada flanco actualiza el estado del controlador)
   SYNC_PROC: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (reset = '1') then
            state <= INI;
         else
            state <= next_state;
         end if;        
      end if;
   end process;
 
--MEALY State-Machine - Outputs based on state and inputs
   OUTPUT_DECODE: process (state) --IMPORTANTE: hay que poner en la lista de sensibilidad todas las se�ales de entrada de este proceso (que es un m�dulo combinacional)
   begin
-- valores por defecto, si no se asigna otro valor en un estado valdr�n lo que se asigna aqu�
		  update_done <= '0';
		  reset_count <= '0';
		  count_enable <= '0';
		  load_data <= '0';
		  DMA_MD_RE <= '0';
		  DMA_MD_WE <= '0';
		  DMA_IO_RE <= '0';
		  DMA_IO_WE <= '0';
		  DMA_sync <= '0';
		  DMA_send_data <= '0';
		  DMA_send_addr <= '0';
		  DMA_Burst <= '0';
		  DMA_wait <= '0';
          next_state <= state;  
        if (state = INI) then -- si no piden nada no hacemos nada
        	
       elsif (state = Escribir_IO) then 
       
       elsif (state = Leer_IO) then 
         	
	   else 
	   end if;
   end process;
 
   
end Behavioral;

